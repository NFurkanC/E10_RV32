`include "../include/rv32_opcodes.vh"

module LSU (
    input wire [:] ,
)