//INCOMPLETE - SUBJECT TO CHANGES
//BARE SKELETON TO FILL FILE STRUCTURE
`include "../include/rv32_opcodes.vh"

module core_control (
    input [31:0] opcode_in,
    output wire regfile_write_en_out,
    
);
    
endmodule