//INCOMPLETE - SUBJECT TO CHANGES
//BARE SKELETON TO FILL FILE STRUCTURE
`include "../include/rv32_opcodes.vh"

module core_top (
    
);

endmodule