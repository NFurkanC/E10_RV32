`ifndef RISCV_32_OPCODES
`define RISCV_32_OPCODES

`define OP_LUI 32'b?????????????????????????0110111
`define OP_AUIPC 32'b?????????????????????????0010111
`define OP_ADDI 32'b?????????????????000?????0010011
`define OP_SLTI 32'b?????????????????010?????0010011
`define OP_SLTIU 32'b?????????????????011?????0010011
`define OP_XORI 32'b?????????????????100?????0010011
`define OP_ORI 32'b?????????????????110?????0010011
`define OP_ANDI 32'b?????????????????111?????0010011
`define OP_SLLI 32'b0000000??????????001?????0010011
`define OP_SRLI 32'b0000000??????????101?????0010011
`define OP_SRAI 32'b0100000??????????101?????0010011
`define OP_ADD 32'b0000000??????????000?????0110011
`define OP_SUB 32'b0100000??????????000?????0110011
`define OP_SLL 32'b0000000??????????001?????0110011
`define OP_SLT 32'b0000000??????????010?????0110011
`define OP_SLTU 32'b0000000??????????011?????0110011
`define OP_XOR 32'b0000000??????????100?????0110011
`define OP_SRL 32'b0000000??????????101?????0110011
`define OP_SRA 32'b0100000??????????101?????0110011
`define OP_OR 32'b0000000??????????110?????0110011
`define OP_AND 32'b0000000??????????111?????0110011
`define OP_FENCE 32'b????????????00000000000000001111
`define OP_FENCE.I 32'b00000000000000000001000000001111
`define OP_CSRRW 32'b?????????????????001?????1110011
`define OP_CSRRS 32'b?????????????????010?????1110011
`define OP_CSRRC 32'b?????????????????011?????1110011
`define OP_CSRRWI 32'b?????????????????101?????1110011
`define OP_CSRRSI 32'b?????????????????110?????1110011
`define OP_CSRRCI 32'b?????????????????111?????1110011
`define OP_ECALL 32'b00000000000000000000000001110011
`define OP_EBREAK 32'b00000000000100000000000001110011
`define OP_URET 0
`define OP_SRET 0
`define OP_MRET 32'b00110000001000000000000001110011
`define OP_WFI 32'b00010000010100000000000001110011
`define OP_SFENCE.VMA
`define OP_LB 32'b?????????????????000?????0000011
`define OP_LH 32'b?????????????????001?????0000011
`define OP_LW 32'b?????????????????010?????0000011
`define OP_LBU 32'b?????????????????100?????0000011
`define OP_LHU 32'b?????????????????101?????0000011
`define OP_SB 32'b?????????????????000?????0100011
`define OP_SH 32'b?????????????????001?????0100011
`define OP_SW 32'b?????????????????010?????0100011
`define OP_JAL 32'b?????????????????????????1101111
`define OP_JALR 32'b?????????????????000?????1100111
`define OP_BEQ 32'b?????????????????000?????1100011
`define OP_BNE 32'b?????????????????001?????1100011
`define OP_BLT 32'b?????????????????100?????1100011
`define OP_BGE 32'b?????????????????101?????1100011
`define OP_BLTU 32'b?????????????????110?????1100011
`define OP_BGEU 32'b?????????????????111?????1100011

//ALU SUBOPCODES

`define ALU_ADD 4'b0000
`define ALU_SUB 4'b0001
`define ALU_AND 4'b0010
`define ALU_OR 4'b0011
`define ALU_XOR 4'b0100
`define ALU_SLL 4'b0101
`define ALU_SRL 4'b0110
`define ALU_SRA 4'b0111
`define ALU_SLT 4'b1000
`define ALU_SLTA 4'b1001

`endif