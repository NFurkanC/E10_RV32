//INCOMPLETE - SUBJECT TO CHANGES
//BARE SKELETON TO FILL FILE STRUCTURE
module top (
  input clk_i,
  input rst_i
);

  wire [31:0] instr;
  wire [31:0] instr_addr;
  wire [31:0] data;
  wire [31:0] data_addr;

endmodule
